//-----------------------------------------------------------------------------
// This program is free software; you can redistribute it and/or
// modify it under the terms of the GNU General Public License
// as published by the Free Software Foundation; either version 2
// of the License, or (at your option) any later version.
//
// This program is distributed in the hope that it will be useful,
// but WITHOUT ANY WARRANTY; without even the implied warranty of
// MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
// GNU General Public License for more details.
//
// You should have received a copy of the GNU General Public License
// along with this program; if not, write to the Free Software
// Foundation, Inc., 51 Franklin Street, Fifth Floor
// Boston, MA  02110-1301, USA.
//
// You can dowload a copy of the GNU General Public License here:
// http://www.gnu.org/licenses/gpl.txt
//
// Copyright (c) March 2022 CERN

//-----------------------------------------------------------------------------
// @file BUILD_NUMBER.SV
// @brief SHOULD BE AUTOGENERATED
// @author Dr. David Belohrad  <david@belohrad.ch>, CERN
// @date 11 March 2022
// @details
// but is not yet for Xilinx
//
// @platform Altera Quartus
// @standard IEEE 1800-2012
//-----------------------------------------------------------------------------

import CKRSPkg::*;


module build_number

  (output logic [31:0] build_ob32
   );

   assign build_ob32 = 32'haabbccdd;





endmodule // build_number
